.SUBCKT INV I ZN
MM1 ZN I VDD VDD pmos_rvt w=162.00n l=20n nfin=6
MM2 ZN I VSS VSS nmos_rvt w=81.0n l=20n nfin=3
.ENDS